--none1
